library IEEE;

use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity project_reti_logiche is
    port (
        i_clk           : in std_logic;
        i_rst           : in std_logic;
        i_start         : in std_logic;
        i_w             : in std_logic;
        o_z0            : out std_logic_vector(7 downto 0);
        o_z1            : out std_logic_vector(7 downto 0);
        o_z2            : out std_logic_vector(7 downto 0);
        o_z3            : out std_logic_vector(7 downto 0);
        o_done          : out std_logic;
        o_mem_addr      : out std_logic_vector(15 downto 0);
        i_mem_data      : in std_logic_vector(7 downto 0);
        o_mem_we        : out std_logic;
        o_mem_en        : out std_logic
    );
end project_reti_logiche;